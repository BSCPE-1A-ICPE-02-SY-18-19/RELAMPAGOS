CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 170 1 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
10
2 +V
167 329 521 0 1 3
0 2
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5130 0 0
2
43530.3 0
0
6 74LS48
188 814 551 0 14 29
0 5 7 9 3 34 35 16 15 14
13 12 11 10 36
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U7
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
391 0 0
2
43530.3 0
0
9 2-In AND~
219 649 504 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3124 0 0
2
43530.3 0
0
9 2-In AND~
219 522 495 0 3 22
0 3 9 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3421 0 0
2
43530.3 0
0
6 74112~
219 714 636 0 7 32
0 2 6 4 6 2 37 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U6B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 5 0
1 U
8157 0 0
2
43530.3 0
0
6 74112~
219 584 635 0 7 32
0 2 8 4 8 2 38 7
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U6A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 5 0
1 U
5572 0 0
2
43530.3 0
0
6 74112~
219 446 635 0 7 32
0 2 3 4 3 2 39 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U5B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 4 0
1 U
8901 0 0
2
43530.3 0
0
6 74112~
219 328 635 0 7 32
0 2 40 4 41 2 42 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U5A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
7361 0 0
2
43530.3 0
0
7 Pulser~
4 250 608 0 10 12
0 43 44 45 4 0 0 5 5 1
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4747 0 0
2
43530.3 0
0
9 CC 7-Seg~
183 898 459 0 18 19
10 29 28 27 26 25 24 23 55 56
1 0 0 1 0 1 1 2 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
972 0 0
2
43530.3 1
0
35
13 1 0 0 0 0 0 2 10 0 0 3
846 569
877 569
877 495
12 2 0 0 0 0 0 2 10 0 0 3
846 560
883 560
883 495
11 3 0 0 0 0 0 2 10 0 0 3
846 551
889 551
889 495
10 4 0 0 0 0 0 2 10 0 0 3
846 542
895 542
895 495
9 5 0 0 0 0 0 2 10 0 0 3
846 533
901 533
901 495
8 6 0 0 0 0 0 2 10 0 0 3
846 524
907 524
907 495
7 7 0 0 0 0 0 2 10 0 0 3
846 515
913 515
913 495
0 0 2 0 0 4096 0 0 0 20 13 2
376 555
376 707
0 0 2 0 0 0 0 0 0 20 12 2
511 555
511 707
0 0 2 0 0 0 0 0 0 20 11 2
668 555
668 707
0 5 2 0 0 0 0 0 5 12 0 3
584 707
714 707
714 648
0 5 2 0 0 0 0 0 6 13 0 3
446 707
584 707
584 647
5 5 2 0 0 16 0 8 7 0 0 4
328 647
328 707
446 707
446 647
0 1 3 0 0 4096 0 0 4 15 0 3
403 617
403 486
498 486
4 2 3 0 0 0 0 7 7 0 0 4
422 617
403 617
403 599
422 599
3 3 4 0 0 12416 0 7 6 0 0 6
416 608
412 608
412 668
546 668
546 608
554 608
1 0 2 0 0 0 0 1 0 0 20 2
329 530
329 555
1 0 2 0 0 0 0 6 0 0 20 2
584 572
584 555
1 0 2 0 0 0 0 7 0 0 20 2
446 572
446 555
1 1 2 0 0 8320 0 5 8 0 0 4
714 573
714 555
328 555
328 572
7 1 5 0 0 8320 0 5 2 0 0 4
738 600
776 600
776 515
782 515
2 3 6 0 0 8320 0 5 3 0 0 4
690 600
684 600
684 504
670 504
2 4 6 0 0 0 0 5 5 0 0 4
690 600
684 600
684 618
690 618
7 2 7 0 0 12416 0 6 2 0 0 4
608 599
658 599
658 524
782 524
7 2 7 0 0 0 0 6 3 0 0 4
608 599
618 599
618 513
625 513
4 2 8 0 0 8192 0 6 6 0 0 4
560 617
555 617
555 599
560 599
2 3 8 0 0 8320 0 6 4 0 0 4
560 599
555 599
555 495
543 495
7 4 3 0 0 12416 0 8 2 0 0 4
352 599
391 599
391 542
782 542
7 3 9 0 0 12416 0 7 2 0 0 4
470 599
540 599
540 533
782 533
7 2 9 0 0 0 0 7 4 0 0 4
470 599
487 599
487 504
498 504
7 2 3 0 0 0 0 8 7 0 0 2
352 599
422 599
3 4 4 0 0 0 0 8 9 0 0 2
298 608
280 608
3 3 4 0 0 0 0 6 5 0 0 6
554 608
550 608
550 668
676 668
676 609
684 609
3 3 4 0 0 0 0 8 7 0 0 6
298 608
294 608
294 668
408 668
408 608
416 608
3 1 8 0 0 0 0 4 3 0 0 2
543 495
625 495
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
349 279 450 303
359 287 439 303
10 Relampagos
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
218 279 367 303
228 287 356 303
16 Joseph Caesar O.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
441 279 526 303
451 287 515 303
8 BSCpE-1A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
